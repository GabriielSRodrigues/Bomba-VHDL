package Common is

  TYPE BombaStage is (armando, contagem, defused, exploded);

end Common;
 
